module toplevel(input CLOCK_50,
					 )

endmodule;